module hi;

initial begin
	$display("hiya");
	#10 $finish;
end

endmodule
